
//--------------------------------------------------------------------------------------------------------
// fpga_top
// Тип     : синтезируемый, верхний уровень FPGA
// Стандарт: Verilog 2001 (IEEE1364-2001)
// Функция : пример использования FOC, верхний модуль проекта FPGA. Управляет тангенциальным моментом двигателя —
//           то по часовой стрелке, то против часовой стрелки. Также можно через UART наблюдать кривую
//           отклика контура тока.
//--------------------------------------------------------------------------------------------------------

module fpga_top (
    input  wire clk_50m, // подключение к кварцевому генератору 50 МГц
    // ------- 3-фазные PWM сигналы (включая сигнал разрешения) ------------------------------------------
    output wire pwm_en,  // общий сигнал разрешения для 3 фаз; если pwm_en=0, все 6 MOSFET закрыты
    output wire pwm_a,   // PWM сигнал фазы A; =0 → открыт нижний транзистор, =1 → открыт верхний транзистор
    output wire pwm_b,   // PWM сигнал фазы B; =0 → открыт нижний транзистор, =1 → открыт верхний транзистор
    output wire pwm_c,   // PWM сигнал фазы C; =0 → открыт нижний транзистор, =1 → открыт верхний транзистор
    // ------- AD7928 (чип АЦП), используется для измерения фазных токов (SPI интерфейс) -----------------
    output wire spi_ss,
    output wire spi_sck,
    output wire spi_mosi,
    input  wire spi_miso,
    // ------- Магнитный энкодер AS5600, используется для получения механического угла ротора (I2C) -------
    output wire i2c_scl,
    inout       i2c_sda,
    // ------- UART: вывод значений реального и целевого тока d-оси (id, id_aim) и q-оси (iq, iq_aim) ----
    output wire uart_tx
);


wire               rstn;        // сигнал сброса, изначально 0; после успешной PLL-синхронизации устанавливается в 1
wire               clk;         // тактовый сигнал (десятки МГц). Частота управления = частота тактирования / 2048.
                                // Например, при 36.864 МГц → частота управления = 36.864МГц/2048 = 18 кГц.
                                // (частота управления = частота дискретизации 3-фазного тока = частота PID-регулятора = частота обновления ШИМ SVPWM)

wire        [11:0] phi;         // механический угол ротора φ, считанный с AS5600, диапазон 0~4095.
                                // 0 → 0°; 1024 → 90°; 2048 → 180°; 3072 → 270°

wire               sn_adc;      // управляющий сигнал момента выборки 3-фазного тока.
                                // Когда требуется выборка, на sn_adc формируется импульс высокого уровня на один такт.
wire               en_adc;      // сигнал готовности результата АЦП.
                                // После импульса sn_adc модуль adc_ad7928 начинает выборку,
                                // по окончании преобразования выдает импульс en_adc и значения токов (adc_value_a/b/c).
wire        [11:0] adc_value_a; // исходное значение АЦП для тока фазы A
wire        [11:0] adc_value_b; // исходное значение АЦП для тока фазы B
wire        [11:0] adc_value_c; // исходное значение АЦП для тока фазы C

wire               en_idq;      // импульс высокого уровня указывает, что появились новые значения id и iq;
                                // каждый цикл управления генерируется один импульс
wire signed [15:0] id;          // фактическое значение тока по d-оси ротора (прямая ось)
wire signed [15:0] iq;          // фактическое значение тока по q-оси ротора (квадратурная ось), может быть положительным или отрицательным
                                // (например: положительное → против часовой стрелки, отрицательное → по часовой, или наоборот)
wire signed [15:0] id_aim;      // целевое значение тока по d-оси, может быть положительным или отрицательным
reg  signed [15:0] iq_aim;      // целевое значение тока по q-оси, может быть положительным или отрицательным
                                // (например: положительное → против часовой стрелки, отрицательное → по часовой, или наоборот)

// PLL использует тактовую частоту 50 МГц (clk_50m) для генерации тактовой частоты 36,864 МГц (clk)
// Примечание: Этот модуль применим только к ПЛИС Altera Cyclone IV. Для ПЛИС других производителей или серий используйте эквивалентные IP-ядра/примитивы (например, Clock Wizard от Xilinx) вместо этого модуля.
wire [3:0] subwire0;
altpll u_altpll ( .inclk ( {1'b0, clk_50m} ), .clk ( {subwire0, clk} ), .locked ( rstn ),  .activeclock (),  .areset (1'b0), .clkbad (),  .clkena ({6{1'b1}}),  .clkloss (), .clkswitch (1'b0), .configupdate (1'b0), .enable0 (), .enable1 (),  .extclk (),  .extclkena ({4{1'b1}}), .fbin (1'b1), .fbmimicbidir (),  .fbout (), .fref (), .icdrclk (), .pfdena (1'b1), .phasecounterselect ({4{1'b1}}), .phasedone (), .phasestep (1'b1), .phaseupdown (1'b1),  .pllena (1'b1), .scanaclr (1'b0), .scanclk (1'b0), .scanclkena (1'b1), .scandata (1'b0), .scandataout (),  .scandone (), .scanread (1'b0), .scanwrite (1'b0), .sclkout0 (), .sclkout1 (), .vcooverrange (), .vcounderrange ());
defparam u_altpll.bandwidth_type = "AUTO", u_altpll.clk0_divide_by = 99,  u_altpll.clk0_duty_cycle = 50, u_altpll.clk0_multiply_by = 73, u_altpll.clk0_phase_shift = "0", u_altpll.compensate_clock = "CLK0", u_altpll.inclk0_input_frequency = 20000, u_altpll.intended_device_family = "Cyclone IV E",  u_altpll.lpm_hint = "CBX_MODULE_PREFIX=pll", u_altpll.lpm_type = "altpll",  u_altpll.operation_mode = "NORMAL",  u_altpll.pll_type = "AUTO", u_altpll.port_activeclock = "PORT_UNUSED",  u_altpll.port_areset = "PORT_UNUSED",  u_altpll.port_clkbad0 = "PORT_UNUSED",  u_altpll.port_clkbad1 = "PORT_UNUSED", u_altpll.port_clkloss = "PORT_UNUSED", u_altpll.port_clkswitch = "PORT_UNUSED", u_altpll.port_configupdate = "PORT_UNUSED", u_altpll.port_fbin = "PORT_UNUSED", u_altpll.port_inclk0 = "PORT_USED",  u_altpll.port_inclk1 = "PORT_UNUSED", u_altpll.port_locked = "PORT_USED", u_altpll.port_pfdena = "PORT_UNUSED",  u_altpll.port_phasecounterselect = "PORT_UNUSED", u_altpll.port_phasedone = "PORT_UNUSED", u_altpll.port_phasestep = "PORT_UNUSED", u_altpll.port_phaseupdown = "PORT_UNUSED",  u_altpll.port_pllena = "PORT_UNUSED", u_altpll.port_scanaclr = "PORT_UNUSED",  u_altpll.port_scanclk = "PORT_UNUSED", u_altpll.port_scanclkena = "PORT_UNUSED", u_altpll.port_scandata = "PORT_UNUSED", u_altpll.port_scandataout = "PORT_UNUSED", u_altpll.port_scandone = "PORT_UNUSED", u_altpll.port_scanread = "PORT_UNUSED", u_altpll.port_scanwrite = "PORT_UNUSED", u_altpll.port_clk0 = "PORT_USED", u_altpll.port_clk1 = "PORT_UNUSED", u_altpll.port_clk2 = "PORT_UNUSED",  u_altpll.port_clk3 = "PORT_UNUSED", u_altpll.port_clk4 = "PORT_UNUSED", u_altpll.port_clk5 = "PORT_UNUSED", u_altpll.port_clkena0 = "PORT_UNUSED",  u_altpll.port_clkena1 = "PORT_UNUSED", u_altpll.port_clkena2 = "PORT_UNUSED", u_altpll.port_clkena3 = "PORT_UNUSED",  u_altpll.port_clkena4 = "PORT_UNUSED", u_altpll.port_clkena5 = "PORT_UNUSED", u_altpll.port_extclk0 = "PORT_UNUSED", u_altpll.port_extclk1 = "PORT_UNUSED",  u_altpll.port_extclk2 = "PORT_UNUSED",  u_altpll.port_extclk3 = "PORT_UNUSED",  u_altpll.self_reset_on_loss_lock = "OFF",  u_altpll.width_clock = 5;
//assign rstn=1'b1; assign clk=clk_50m;


// Простой контроллер чтения I2C, реализует чтение магнитного энкодера AS5600, считывает текущий механический угол ротора φ
wire [3:0] i2c_trash;    // отбрасываем старшие 4 бита
i2c_register_read #(
    .CLK_DIV      ( 16'd10         ),  // коэффициент деления тактового сигнала i2c_scl, частота scl = частота clk / (4*CLK_DIV). Например, в этом примере clk равен 36,864 МГц, CLK_DIV = 10, тогда частота SCL равна 36864/(4*10) = 922 кГц. Примечание: для микросхемы AS5600 требуется частота SCL не более 1 МГц.
    .SLAVE_ADDR   ( 7'h36          ),  // AS5600's I2C slave address
    .REGISTER_ADDR( 8'h0E          )   // the register address to read
) u_as5600_read (
    .rstn         ( rstn           ),
    .clk          ( clk            ),
    .scl          ( i2c_scl        ), // Интерфейс I2C: SCL
    .sda          ( i2c_sda        ), // Интерфейс I2C: SDA
    .start        ( 1'b1           ), // Продолжить операцию чтения I2C
    .ready        (                ),
    .done         (                ),
    .regout       ( {i2c_trash, phi} )
);



// Считыватель АЦП AD7928, используемый для считывания значений выборки трёхфазного тока (необработанные значения АЦП считываются без какой-либо обработки)
adc_ad7928 #(
    .CH_CNT       ( 3'd2           ), // Этот параметр установлен в 2, что указывает на то, что нам нужны только значения АЦП CH0, CH1 и CH2
    .CH0          ( 3'd1           ), // Указывает, что CH0 соответствует каналу 1 AD7928. (Аппаратно ток фазы A подключен к каналу 1 AD7928)
    .CH1          ( 3'd2           ), // Указывает, что CH1 соответствует каналу 2 AD7928. (Аппаратно ток фазы B подключен к каналу 2 AD7928)
    .CH2          ( 3'd3           )  // Указывает, что CH2 соответствует каналу 3 AD7928. (Аппаратно ток фазы C подключен к AD7928 канал 3)
) u_adc_ad7928 (
    .rstn         ( rstn           ),
    .clk          ( clk            ),
    .spi_ss       ( spi_ss         ), // Интерфейс SPI: SS
    .spi_sck      ( spi_sck        ), // Интерфейс SPI: SCK
    .spi_mosi     ( spi_mosi       ), // Интерфейс SPI: MOSI
    .spi_miso     ( spi_miso       ), // Интерфейс SPI: MISO
    .i_sn_adc     ( sn_adc         ), // input : Когда sn_adc формирует импульс высокого уровня, модуль начинает (трёхканальное) преобразование АЦП
    .o_en_adc     ( en_adc         ), // output: После завершения преобразования en_adc формирует период импульсов высокого уровня
    .o_adc_value0 ( adc_value_a    ), // Когда en_adc формирует период высокоуровневых импульсов, adc_value_a отображается как необработанное значение АЦП фазных токов
    .o_adc_value1 ( adc_value_b    ), // Когда en_adc формирует высокоуровневый импульс в течение одного цикла, необработанное значение АЦП тока фазы B отображается на adc_value_b
    .o_adc_value2 ( adc_value_c    ), // Когда en_adc формирует высокоуровневый импульс в течение одного цикла, необработанное значение АЦП тока фазы C отображается на adc_value_c
    .o_adc_value3 (                ), // Игнорируем оставшиеся пять результатов преобразования АЦП
    .o_adc_value4 (                ), // Игнорируем оставшиеся пять результатов преобразования АЦП
    .o_adc_value5 (                ), // Игнорируем оставшиеся пять результатов преобразования АЦП
    .o_adc_value6 (                ), // Игнорируем оставшиеся пять результатов преобразования АЦП
    .o_adc_value7 (                )  // Игнорируем оставшиеся пять результатов преобразования АЦП
);



// Модуль FOC + SVPWM (Подробное использование и принципы работы см. в файле foc_top.sv)
foc_top #(
    .INIT_CYCLES  ( 16777216       ), // В этом примере тактовая частота (clk) составляет 36,864 МГц. Если INIT_CYCLES = 16777216, время инициализации составляет 16777216/36864000 = 0,45 секунды.
    .ANGLE_INV    ( 1'b0           ), // В этом примере датчик угла установлен не в перевёрнутом виде (направление вращения A->B->C->A совпадает с направлением увеличения φ), поэтому этот параметр следует установить равным 0.
    .POLE_PAIR    ( 8'd7           ), // Количество пар полюсов, используемых в этом примере, равно 7.
    .MAX_AMP      ( 9'd384         ), // 384 / 512 = 0,75. Это означает, что максимальная амплитуда SVPWM составляет 75% от максимального предела амплитуды.
    .SAMPLE_DELAY ( 9'd120         )  // Задержка выборки, диапазон значений 0–511. Учитывая, что трёхфазным МОП-транзисторам драйверам требуется время для стабилизации после начала включения тока, требуется определённая задержка между моментом включения всех трёх нижних плеч моста и моментом выборки АЦП. Этот параметр определяет количество тактовых циклов этой задержки. По окончании задержки модуль формирует импульс высокого уровня на сигнале sn_adc, указывая на готовность внешнего АЦП к выборке.
) u_foc_top (
    .rstn         ( rstn           ),
    .clk          ( clk            ),
    .Kp           ( 31'd300000     ), // Параметр P для алгоритма ПИД-регулирования токового контура
    .Ki           ( 31'd30000      ), // Параметр I для ПИД-регулирования токового контура Алгоритма
    .phi          ( phi            ), // input: Вход датчика угла (механический угол, сокращённо φ), диапазон значений от 0 до 4095. 0 соответствует 0°; 1024 соответствует 90°; 2048 соответствует 180°; а 3072 соответствует 270°.
    .sn_adc       ( sn_adc         ), // output: Сигнал управления тактовой частотой дискретизации трёхфазного АЦП тока. При необходимости выборки на сигнале sn_adc формируется импульс высокого уровня длительностью в один такт, указывая на необходимость начала выборки АЦП.
    .en_adc       ( en_adc         ), // input : Сигнал подтверждения результата выборки трёхфазного АЦП тока. После формирования импульса высокого уровня на сигнале sn_adc внешний АЦП начинает выборку трёхфазного тока. После завершения преобразования на сигнале en_adc должен быть сформирован импульс высокого уровня длительностью в один такт. Одновременно с этим выполняется преобразование АЦП. Результат формируется на основе сигналов adc_a, adc_b и adc_c.
    .adc_a        ( adc_value_a    ), // input : Результат выборки АЦП фазы A
    .adc_b        ( adc_value_b    ), // input : Результат выборки АЦП фазы B
    .adc_c        ( adc_value_c    ), // input : Результат выборки АЦП фазы C
    .pwm_en       ( pwm_en         ),
    .pwm_a        ( pwm_a          ),
    .pwm_b        ( pwm_b          ),
    .pwm_c        ( pwm_c          ),
    .en_idq       ( en_idq         ), // output: Импульс высокого уровня указывает на то, что id и iq получили новые значения. en_idq генерирует импульс высокого уровня в течение каждого цикла управления
    .id           ( id             ), // output: d Фактическое значение тока по оси d (ось ординат), может быть положительным или отрицательным
    .iq           ( iq             ), // output: q Фактическое значение тока по оси q (квадратурной оси), может быть положительным или отрицательным (положительное значение соответствует вращению против часовой стрелки, отрицательное — по часовой стрелке, и наоборот).
    .id_aim       ( id_aim         ), // input : d Целевое значение тока по оси d (прямой оси), может быть положительным или отрицательным. Обычно устанавливается равным 0, если управление ослаблением поля не используется.
    .iq_aim       ( iq_aim         ), // input : q Целевое значение тока по оси q (прямой оси), может быть положительным или отрицательным (положительное значение соответствует вращению против часовой стрелки, отрицательное — по часовой стрелке, и наоборот).
    .init_done    (                )  // output: Сигнал завершения инициализации. До завершения инициализации = 0; после завершения инициализации (переход в состояние управления FOC) = 1
);



reg [23:0] cnt;
always @ (posedge clk or negedge rstn)   // Этот always-блок реализует 24-битный счётчик с автоинкрементом
    if(~rstn)
        cnt <= 24'd0;
    else
        cnt <= cnt + 24'd1;


assign id_aim = $signed(16'd0);          // Задаём id_aim равным 0 постоянно

always @ (posedge clk or negedge rstn)   // Этот always-блок попеременно присваивает iq_aim значения +200 и -200,
    if(~rstn) begin                      // то есть тангенциальный момент двигателя меняется то по часовой стрелке, то против часовой
        iq_aim <= $signed(16'd0);
    end else begin
        if(cnt[23])
            iq_aim <=  $signed(16'd200); // 令 id_aim = +200
        else
            iq_aim <= -$signed(16'd200); // 令 id_aim = -200
    end



// UART передатчик (монитор), формат: 115200,8,n,1
uart_monitor #(
    .CLK_DIV      ( 16'd320        )   // коэффициент деления UART, здесь 320.
                                        // Так как частота тактового сигнала 36.864 МГц, то 36.864МГц / 320 = 115200 бод
) u_uart_monitor (
    .rstn         ( rstn           ),
    .clk          ( clk            ),
    .i_en         ( en_idq         ),  // input: при появлении импульса высокого уровня на en_idq запускается передача по UART
    .i_val0       ( id             ),  // input: отправка переменной id в десятичном виде
    .i_val1       ( id_aim         ),  // input: отправка переменной id_aim в десятичном виде
    .i_val2       ( iq             ),  // input: отправка переменной iq в десятичном виде
    .i_val3       ( iq_aim         ),  // input: отправка переменной iq_aim в десятичном виде
    .o_uart_tx    ( uart_tx        )   // output: выходной сигнал UART передачи
);


endmodule
